LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY DE2LAB1 IS
	PORT(
		SW : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
		HEX0: OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
		HEX1: OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
		HEX2: OUT STD_LOGIC_VECTOR(6 DOWNTO 0)
	);
END ENTITY;

ARCHITECTURE STRUCT OF DE2LAB1 IS
--COMPONENT DECLARATION
COMPONENT DECODER IS
	PORT(
		SW : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
		MUX : OUT STD_LOGIC_VECTOR(5 DOWNTO 0)
	);
END COMPONENT;

COMPONENT MUX IS
	PORT(
		SW0 : IN STD_LOGIC_VECTOR(9 DOWNTO 8);
		SW1 : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		MUX0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0)
	);
END COMPONENT;

COMPONENT SEGMENT7 IS
	PORT(
		SW : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
		HEX0 : OUT STD_LOGIC_VECTOR(6 DOWNTO 0)
	);
END COMPONENT;

--SIGNAL DECLARATION
SIGNAL DECODED : STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL MUX_0, MUX_1, MUX_2 : STD_LOGIC_VECTOR(1 DOWNTO 0);

BEGIN
	DECODER0 : DECODER PORT MAP( SW(9 DOWNTO 8), DECODED);
	MUX0 : MUX PORT MAP(DECODED(5 DOWNTO 4), SW(5 DOWNTO 0), MUX_0);
	MUX1 : MUX PORT MAP(DECODED(3 DOWNTO 2), SW(5 DOWNTO 0), MUX_1);
	MUX2 : MUX PORT MAP(DECODED(1 DOWNTO 0), SW(5 DOWNTO 0), MUX_2);
	SEG0 : SEGMENT7 PORT MAP(MUX_0, HEX0);
	SEG1 : SEGMENT7 PORT MAP(MUX_1, HEX1);
	SEG2 : SEGMENT7 PORT MAP(MUX_2, HEX2);
END;
