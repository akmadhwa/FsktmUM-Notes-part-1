LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY MUX IS
	PORT(
		SW0: IN STD_LOGIC_VECTOR(9 DOWNTO 8);
		SW1 : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		MUX0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0)
	);
END ENTITY;

ARCHITECTURE STRUCT OF MUX IS	
BEGIN
	PROCESS(SW0,SW1)
	BEGIN	
		IF(SW0(9 DOWNTO 8) = "00")	THEN
			MUX0 <= SW1(5 DOWNTO 4);
		ELSIF(SW0(9 DOWNTO 8) = "01")	THEN
			MUX0 <= SW1(3 DOWNTO 2);
		ELSIF(SW0(9 DOWNTO 8) = "10")	THEN
			MUX0 <= SW1(1 DOWNTO 0);
		END IF;
	END PROCESS;
END ARCHITECTURE STRUCT;