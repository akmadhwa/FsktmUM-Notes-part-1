LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY DECODER IS
	PORT(
		SW : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
		MUX : OUT STD_LOGIC_VECTOR(5 DOWNTO 0)
	);
END ENTITY;

ARCHITECTURE STRUCT OF DECODER IS	
BEGIN
	PROCESS(SW)
	BEGIN
		CASE SW IS
			WHEN "00" => MUX <= "000110";
			WHEN "01" => MUX <= "011000";
			WHEN "10" => MUX <= "100001";
			WHEN "11" => MUX <= "111111";
		END CASE;
	END PROCESS;
END ARCHITECTURE STRUCT;