PACKAGE vm_pack2 IS
	TYPE t_vm_state IS (
		st_r,
		st_g,
		st_y
  
  );
END vm_pack;