LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY SEGMENT7 IS
	PORT(
		SW : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
		HEX0 : OUT STD_LOGIC_VECTOR(6 DOWNTO 0)
	);
END ENTITY;

ARCHITECTURE STRUCT OF SEGMENT7 IS	
BEGIN
	PROCESS(SW)
	BEGIN
		CASE SW IS
			WHEN "00" => HEX0 <= "0100001";
			WHEN "01" => HEX0 <= "0000110";
			WHEN "10" => HEX0 <= "0100100";
			WHEN "11" => HEX0 <= "1111111";
		END CASE;
	END PROCESS;
END ARCHITECTURE STRUCT;